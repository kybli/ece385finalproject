module audio_mux (	input logic [10:0] AVL_ADDR,
					input logic [31:0] AVL_WRITEDATA,
					input logic [8191:0] reg_out_packed,
					input logic [31:0] READY_out,
					output logic [31:0] AVL_READDATA,
					output logic READY_load,
					output logic [255:0] fft_load);
always_comb begin
fft_load = 256'b0;
AVL_READDATA = 32'hFFFF;

	case (AVL_ADDR)
		// 10'd0: AVL_READDATA = reg_out_packed[8191 : 8160];
		10'd0: AVL_READDATA = 32'hFFFF;
		// 10'd1: AVL_READDATA = reg_out_packed[8159 : 8128];
		10'd1: AVL_READDATA = 32'hFFFF;
		// 10'd2: AVL_READDATA = reg_out_packed[8127 : 8096];
		10'd2: AVL_READDATA = 32'hFFFF;
		// 10'd3: AVL_READDATA = reg_out_packed[8095 : 8064];
		10'd3: AVL_READDATA = 32'hFFFF;
		10'd4: AVL_READDATA = reg_out_packed[8063 : 8032];
		10'd5: AVL_READDATA = reg_out_packed[8031 : 8000];
		10'd6: AVL_READDATA = reg_out_packed[7999 : 7968];
		10'd7: AVL_READDATA = reg_out_packed[7967 : 7936];
		10'd8: AVL_READDATA = reg_out_packed[7935 : 7904];
		10'd9: AVL_READDATA = reg_out_packed[7903 : 7872];
		10'd10: AVL_READDATA = reg_out_packed[7871 : 7840];
		10'd11: AVL_READDATA = reg_out_packed[7839 : 7808];
		10'd12: AVL_READDATA = reg_out_packed[7807 : 7776];
		10'd13: AVL_READDATA = reg_out_packed[7775 : 7744];
		10'd14: AVL_READDATA = reg_out_packed[7743 : 7712];
		10'd15: AVL_READDATA = reg_out_packed[7711 : 7680];
		10'd16: AVL_READDATA = reg_out_packed[7679 : 7648];
		10'd17: AVL_READDATA = reg_out_packed[7647 : 7616];
		10'd18: AVL_READDATA = reg_out_packed[7615 : 7584];
		10'd19: AVL_READDATA = reg_out_packed[7583 : 7552];
		10'd20: AVL_READDATA = reg_out_packed[7551 : 7520];
		10'd21: AVL_READDATA = reg_out_packed[7519 : 7488];
		10'd22: AVL_READDATA = reg_out_packed[7487 : 7456];
		10'd23: AVL_READDATA = reg_out_packed[7455 : 7424];
		10'd24: AVL_READDATA = reg_out_packed[7423 : 7392];
		10'd25: AVL_READDATA = reg_out_packed[7391 : 7360];
		10'd26: AVL_READDATA = reg_out_packed[7359 : 7328];
		10'd27: AVL_READDATA = reg_out_packed[7327 : 7296];
		10'd28: AVL_READDATA = reg_out_packed[7295 : 7264];
		10'd29: AVL_READDATA = reg_out_packed[7263 : 7232];
		10'd30: AVL_READDATA = reg_out_packed[7231 : 7200];
		10'd31: AVL_READDATA = reg_out_packed[7199 : 7168];
		10'd32: AVL_READDATA = reg_out_packed[7167 : 7136];
		10'd33: AVL_READDATA = reg_out_packed[7135 : 7104];
		10'd34: AVL_READDATA = reg_out_packed[7103 : 7072];
		10'd35: AVL_READDATA = reg_out_packed[7071 : 7040];
		10'd36: AVL_READDATA = reg_out_packed[7039 : 7008];
		10'd37: AVL_READDATA = reg_out_packed[7007 : 6976];
		10'd38: AVL_READDATA = reg_out_packed[6975 : 6944];
		10'd39: AVL_READDATA = reg_out_packed[6943 : 6912];
		10'd40: AVL_READDATA = reg_out_packed[6911 : 6880];
		10'd41: AVL_READDATA = reg_out_packed[6879 : 6848];
		10'd42: AVL_READDATA = reg_out_packed[6847 : 6816];
		10'd43: AVL_READDATA = reg_out_packed[6815 : 6784];
		10'd44: AVL_READDATA = reg_out_packed[6783 : 6752];
		10'd45: AVL_READDATA = reg_out_packed[6751 : 6720];
		10'd46: AVL_READDATA = reg_out_packed[6719 : 6688];
		10'd47: AVL_READDATA = reg_out_packed[6687 : 6656];
		10'd48: AVL_READDATA = reg_out_packed[6655 : 6624];
		10'd49: AVL_READDATA = reg_out_packed[6623 : 6592];
		10'd50: AVL_READDATA = reg_out_packed[6591 : 6560];
		10'd51: AVL_READDATA = reg_out_packed[6559 : 6528];
		10'd52: AVL_READDATA = reg_out_packed[6527 : 6496];
		10'd53: AVL_READDATA = reg_out_packed[6495 : 6464];
		10'd54: AVL_READDATA = reg_out_packed[6463 : 6432];
		10'd55: AVL_READDATA = reg_out_packed[6431 : 6400];
		10'd56: AVL_READDATA = reg_out_packed[6399 : 6368];
		10'd57: AVL_READDATA = reg_out_packed[6367 : 6336];
		10'd58: AVL_READDATA = reg_out_packed[6335 : 6304];
		10'd59: AVL_READDATA = reg_out_packed[6303 : 6272];
		10'd60: AVL_READDATA = reg_out_packed[6271 : 6240];
		10'd61: AVL_READDATA = reg_out_packed[6239 : 6208];
		10'd62: AVL_READDATA = reg_out_packed[6207 : 6176];
		10'd63: AVL_READDATA = reg_out_packed[6175 : 6144];
		10'd64: AVL_READDATA = reg_out_packed[6143 : 6112];
		10'd65: AVL_READDATA = reg_out_packed[6111 : 6080];
		10'd66: AVL_READDATA = reg_out_packed[6079 : 6048];
		10'd67: AVL_READDATA = reg_out_packed[6047 : 6016];
		10'd68: AVL_READDATA = reg_out_packed[6015 : 5984];
		10'd69: AVL_READDATA = reg_out_packed[5983 : 5952];
		10'd70: AVL_READDATA = reg_out_packed[5951 : 5920];
		10'd71: AVL_READDATA = reg_out_packed[5919 : 5888];
		10'd72: AVL_READDATA = reg_out_packed[5887 : 5856];
		10'd73: AVL_READDATA = reg_out_packed[5855 : 5824];
		10'd74: AVL_READDATA = reg_out_packed[5823 : 5792];
		10'd75: AVL_READDATA = reg_out_packed[5791 : 5760];
		10'd76: AVL_READDATA = reg_out_packed[5759 : 5728];
		10'd77: AVL_READDATA = reg_out_packed[5727 : 5696];
		10'd78: AVL_READDATA = reg_out_packed[5695 : 5664];
		10'd79: AVL_READDATA = reg_out_packed[5663 : 5632];
		10'd80: AVL_READDATA = reg_out_packed[5631 : 5600];
		10'd81: AVL_READDATA = reg_out_packed[5599 : 5568];
		10'd82: AVL_READDATA = reg_out_packed[5567 : 5536];
		10'd83: AVL_READDATA = reg_out_packed[5535 : 5504];
		10'd84: AVL_READDATA = reg_out_packed[5503 : 5472];
		10'd85: AVL_READDATA = reg_out_packed[5471 : 5440];
		10'd86: AVL_READDATA = reg_out_packed[5439 : 5408];
		10'd87: AVL_READDATA = reg_out_packed[5407 : 5376];
		10'd88: AVL_READDATA = reg_out_packed[5375 : 5344];
		10'd89: AVL_READDATA = reg_out_packed[5343 : 5312];
		10'd90: AVL_READDATA = reg_out_packed[5311 : 5280];
		10'd91: AVL_READDATA = reg_out_packed[5279 : 5248];
		10'd92: AVL_READDATA = reg_out_packed[5247 : 5216];
		10'd93: AVL_READDATA = reg_out_packed[5215 : 5184];
		10'd94: AVL_READDATA = reg_out_packed[5183 : 5152];
		10'd95: AVL_READDATA = reg_out_packed[5151 : 5120];
		10'd96: AVL_READDATA = reg_out_packed[5119 : 5088];
		10'd97: AVL_READDATA = reg_out_packed[5087 : 5056];
		10'd98: AVL_READDATA = reg_out_packed[5055 : 5024];
		10'd99: AVL_READDATA = reg_out_packed[5023 : 4992];
		10'd100: AVL_READDATA = reg_out_packed[4991 : 4960];
		10'd101: AVL_READDATA = reg_out_packed[4959 : 4928];
		10'd102: AVL_READDATA = reg_out_packed[4927 : 4896];
		10'd103: AVL_READDATA = reg_out_packed[4895 : 4864];
		10'd104: AVL_READDATA = reg_out_packed[4863 : 4832];
		10'd105: AVL_READDATA = reg_out_packed[4831 : 4800];
		10'd106: AVL_READDATA = reg_out_packed[4799 : 4768];
		10'd107: AVL_READDATA = reg_out_packed[4767 : 4736];
		10'd108: AVL_READDATA = reg_out_packed[4735 : 4704];
		10'd109: AVL_READDATA = reg_out_packed[4703 : 4672];
		10'd110: AVL_READDATA = reg_out_packed[4671 : 4640];
		10'd111: AVL_READDATA = reg_out_packed[4639 : 4608];
		10'd112: AVL_READDATA = reg_out_packed[4607 : 4576];
		10'd113: AVL_READDATA = reg_out_packed[4575 : 4544];
		10'd114: AVL_READDATA = reg_out_packed[4543 : 4512];
		10'd115: AVL_READDATA = reg_out_packed[4511 : 4480];
		10'd116: AVL_READDATA = reg_out_packed[4479 : 4448];
		10'd117: AVL_READDATA = reg_out_packed[4447 : 4416];
		10'd118: AVL_READDATA = reg_out_packed[4415 : 4384];
		10'd119: AVL_READDATA = reg_out_packed[4383 : 4352];
		10'd120: AVL_READDATA = reg_out_packed[4351 : 4320];
		10'd121: AVL_READDATA = reg_out_packed[4319 : 4288];
		10'd122: AVL_READDATA = reg_out_packed[4287 : 4256];
		10'd123: AVL_READDATA = reg_out_packed[4255 : 4224];
		10'd124: AVL_READDATA = reg_out_packed[4223 : 4192];
		10'd125: AVL_READDATA = reg_out_packed[4191 : 4160];
		10'd126: AVL_READDATA = reg_out_packed[4159 : 4128];
		10'd127: AVL_READDATA = reg_out_packed[4127 : 4096];
		10'd128: AVL_READDATA = reg_out_packed[4095 : 4064];
		10'd129: AVL_READDATA = reg_out_packed[4063 : 4032];
		10'd130: AVL_READDATA = reg_out_packed[4031 : 4000];
		10'd131: AVL_READDATA = reg_out_packed[3999 : 3968];
		10'd132: AVL_READDATA = reg_out_packed[3967 : 3936];
		10'd133: AVL_READDATA = reg_out_packed[3935 : 3904];
		10'd134: AVL_READDATA = reg_out_packed[3903 : 3872];
		10'd135: AVL_READDATA = reg_out_packed[3871 : 3840];
		10'd136: AVL_READDATA = reg_out_packed[3839 : 3808];
		10'd137: AVL_READDATA = reg_out_packed[3807 : 3776];
		10'd138: AVL_READDATA = reg_out_packed[3775 : 3744];
		10'd139: AVL_READDATA = reg_out_packed[3743 : 3712];
		10'd140: AVL_READDATA = reg_out_packed[3711 : 3680];
		10'd141: AVL_READDATA = reg_out_packed[3679 : 3648];
		10'd142: AVL_READDATA = reg_out_packed[3647 : 3616];
		10'd143: AVL_READDATA = reg_out_packed[3615 : 3584];
		10'd144: AVL_READDATA = reg_out_packed[3583 : 3552];
		10'd145: AVL_READDATA = reg_out_packed[3551 : 3520];
		10'd146: AVL_READDATA = reg_out_packed[3519 : 3488];
		10'd147: AVL_READDATA = reg_out_packed[3487 : 3456];
		10'd148: AVL_READDATA = reg_out_packed[3455 : 3424];
		10'd149: AVL_READDATA = reg_out_packed[3423 : 3392];
		10'd150: AVL_READDATA = reg_out_packed[3391 : 3360];
		10'd151: AVL_READDATA = reg_out_packed[3359 : 3328];
		10'd152: AVL_READDATA = reg_out_packed[3327 : 3296];
		10'd153: AVL_READDATA = reg_out_packed[3295 : 3264];
		10'd154: AVL_READDATA = reg_out_packed[3263 : 3232];
		10'd155: AVL_READDATA = reg_out_packed[3231 : 3200];
		10'd156: AVL_READDATA = reg_out_packed[3199 : 3168];
		10'd157: AVL_READDATA = reg_out_packed[3167 : 3136];
		10'd158: AVL_READDATA = reg_out_packed[3135 : 3104];
		10'd159: AVL_READDATA = reg_out_packed[3103 : 3072];
		10'd160: AVL_READDATA = reg_out_packed[3071 : 3040];
		10'd161: AVL_READDATA = reg_out_packed[3039 : 3008];
		10'd162: AVL_READDATA = reg_out_packed[3007 : 2976];
		10'd163: AVL_READDATA = reg_out_packed[2975 : 2944];
		10'd164: AVL_READDATA = reg_out_packed[2943 : 2912];
		10'd165: AVL_READDATA = reg_out_packed[2911 : 2880];
		10'd166: AVL_READDATA = reg_out_packed[2879 : 2848];
		10'd167: AVL_READDATA = reg_out_packed[2847 : 2816];
		10'd168: AVL_READDATA = reg_out_packed[2815 : 2784];
		10'd169: AVL_READDATA = reg_out_packed[2783 : 2752];
		10'd170: AVL_READDATA = reg_out_packed[2751 : 2720];
		10'd171: AVL_READDATA = reg_out_packed[2719 : 2688];
		10'd172: AVL_READDATA = reg_out_packed[2687 : 2656];
		10'd173: AVL_READDATA = reg_out_packed[2655 : 2624];
		10'd174: AVL_READDATA = reg_out_packed[2623 : 2592];
		10'd175: AVL_READDATA = reg_out_packed[2591 : 2560];
		10'd176: AVL_READDATA = reg_out_packed[2559 : 2528];
		10'd177: AVL_READDATA = reg_out_packed[2527 : 2496];
		10'd178: AVL_READDATA = reg_out_packed[2495 : 2464];
		10'd179: AVL_READDATA = reg_out_packed[2463 : 2432];
		10'd180: AVL_READDATA = reg_out_packed[2431 : 2400];
		10'd181: AVL_READDATA = reg_out_packed[2399 : 2368];
		10'd182: AVL_READDATA = reg_out_packed[2367 : 2336];
		10'd183: AVL_READDATA = reg_out_packed[2335 : 2304];
		10'd184: AVL_READDATA = reg_out_packed[2303 : 2272];
		10'd185: AVL_READDATA = reg_out_packed[2271 : 2240];
		10'd186: AVL_READDATA = reg_out_packed[2239 : 2208];
		10'd187: AVL_READDATA = reg_out_packed[2207 : 2176];
		10'd188: AVL_READDATA = reg_out_packed[2175 : 2144];
		10'd189: AVL_READDATA = reg_out_packed[2143 : 2112];
		10'd190: AVL_READDATA = reg_out_packed[2111 : 2080];
		10'd191: AVL_READDATA = reg_out_packed[2079 : 2048];
		10'd192: AVL_READDATA = reg_out_packed[2047 : 2016];
		10'd193: AVL_READDATA = reg_out_packed[2015 : 1984];
		10'd194: AVL_READDATA = reg_out_packed[1983 : 1952];
		10'd195: AVL_READDATA = reg_out_packed[1951 : 1920];
		10'd196: AVL_READDATA = reg_out_packed[1919 : 1888];
		10'd197: AVL_READDATA = reg_out_packed[1887 : 1856];
		10'd198: AVL_READDATA = reg_out_packed[1855 : 1824];
		10'd199: AVL_READDATA = reg_out_packed[1823 : 1792];
		10'd200: AVL_READDATA = reg_out_packed[1791 : 1760];
		10'd201: AVL_READDATA = reg_out_packed[1759 : 1728];
		10'd202: AVL_READDATA = reg_out_packed[1727 : 1696];
		10'd203: AVL_READDATA = reg_out_packed[1695 : 1664];
		10'd204: AVL_READDATA = reg_out_packed[1663 : 1632];
		10'd205: AVL_READDATA = reg_out_packed[1631 : 1600];
		10'd206: AVL_READDATA = reg_out_packed[1599 : 1568];
		10'd207: AVL_READDATA = reg_out_packed[1567 : 1536];
		10'd208: AVL_READDATA = reg_out_packed[1535 : 1504];
		10'd209: AVL_READDATA = reg_out_packed[1503 : 1472];
		10'd210: AVL_READDATA = reg_out_packed[1471 : 1440];
		10'd211: AVL_READDATA = reg_out_packed[1439 : 1408];
		10'd212: AVL_READDATA = reg_out_packed[1407 : 1376];
		10'd213: AVL_READDATA = reg_out_packed[1375 : 1344];
		10'd214: AVL_READDATA = reg_out_packed[1343 : 1312];
		10'd215: AVL_READDATA = reg_out_packed[1311 : 1280];
		10'd216: AVL_READDATA = reg_out_packed[1279 : 1248];
		10'd217: AVL_READDATA = reg_out_packed[1247 : 1216];
		10'd218: AVL_READDATA = reg_out_packed[1215 : 1184];
		10'd219: AVL_READDATA = reg_out_packed[1183 : 1152];
		10'd220: AVL_READDATA = reg_out_packed[1151 : 1120];
		10'd221: AVL_READDATA = reg_out_packed[1119 : 1088];
		10'd222: AVL_READDATA = reg_out_packed[1087 : 1056];
		10'd223: AVL_READDATA = reg_out_packed[1055 : 1024];
		10'd224: AVL_READDATA = reg_out_packed[1023 : 992];
		10'd225: AVL_READDATA = reg_out_packed[991 : 960];
		10'd226: AVL_READDATA = reg_out_packed[959 : 928];
		10'd227: AVL_READDATA = reg_out_packed[927 : 896];
		10'd228: AVL_READDATA = reg_out_packed[895 : 864];
		10'd229: AVL_READDATA = reg_out_packed[863 : 832];
		10'd230: AVL_READDATA = reg_out_packed[831 : 800];
		10'd231: AVL_READDATA = reg_out_packed[799 : 768];
		10'd232: AVL_READDATA = reg_out_packed[767 : 736];
		10'd233: AVL_READDATA = reg_out_packed[735 : 704];
		10'd234: AVL_READDATA = reg_out_packed[703 : 672];
		10'd235: AVL_READDATA = reg_out_packed[671 : 640];
		10'd236: AVL_READDATA = reg_out_packed[639 : 608];
		10'd237: AVL_READDATA = reg_out_packed[607 : 576];
		10'd238: AVL_READDATA = reg_out_packed[575 : 544];
		10'd239: AVL_READDATA = reg_out_packed[543 : 512];
		10'd240: AVL_READDATA = reg_out_packed[511 : 480];
		10'd241: AVL_READDATA = reg_out_packed[479 : 448];
		10'd242: AVL_READDATA = reg_out_packed[447 : 416];
		10'd243: AVL_READDATA = reg_out_packed[415 : 384];
		10'd244: AVL_READDATA = reg_out_packed[383 : 352];
		10'd245: AVL_READDATA = reg_out_packed[351 : 320];
		10'd246: AVL_READDATA = reg_out_packed[319 : 288];
		10'd247: AVL_READDATA = reg_out_packed[287 : 256];
		10'd248: AVL_READDATA = reg_out_packed[255 : 224];
		10'd249: AVL_READDATA = reg_out_packed[223 : 192];
		10'd250: AVL_READDATA = reg_out_packed[191 : 160];
		10'd251: AVL_READDATA = reg_out_packed[159 : 128];
		10'd252: AVL_READDATA = reg_out_packed[127 : 96];
		10'd253: AVL_READDATA = reg_out_packed[95 : 64];
		10'd254: AVL_READDATA = reg_out_packed[63 : 32];
		10'd255: AVL_READDATA = reg_out_packed[31 : 0];
		10'd512: AVL_READDATA = READY_out;
		default: ;
	endcase
	case (AVL_ADDR)
		10'd256: fft_load[0] = 1'b1;
		10'd257: fft_load[1] = 1'b1;
		10'd258: fft_load[2] = 1'b1;
		10'd259: fft_load[3] = 1'b1;
		10'd260: fft_load[4] = 1'b1;
		10'd261: fft_load[5] = 1'b1;
		10'd262: fft_load[6] = 1'b1;
		10'd263: fft_load[7] = 1'b1;
		10'd264: fft_load[8] = 1'b1;
		10'd265: fft_load[9] = 1'b1;
		10'd266: fft_load[10] = 1'b1;
		10'd267: fft_load[11] = 1'b1;
		10'd268: fft_load[12] = 1'b1;
		10'd269: fft_load[13] = 1'b1;
		10'd270: fft_load[14] = 1'b1;
		10'd271: fft_load[15] = 1'b1;
		10'd272: fft_load[16] = 1'b1;
		10'd273: fft_load[17] = 1'b1;
		10'd274: fft_load[18] = 1'b1;
		10'd275: fft_load[19] = 1'b1;
		10'd276: fft_load[20] = 1'b1;
		10'd277: fft_load[21] = 1'b1;
		10'd278: fft_load[22] = 1'b1;
		10'd279: fft_load[23] = 1'b1;
		10'd280: fft_load[24] = 1'b1;
		10'd281: fft_load[25] = 1'b1;
		10'd282: fft_load[26] = 1'b1;
		10'd283: fft_load[27] = 1'b1;
		10'd284: fft_load[28] = 1'b1;
		10'd285: fft_load[29] = 1'b1;
		10'd286: fft_load[30] = 1'b1;
		10'd287: fft_load[31] = 1'b1;
		10'd288: fft_load[32] = 1'b1;
		10'd289: fft_load[33] = 1'b1;
		10'd290: fft_load[34] = 1'b1;
		10'd291: fft_load[35] = 1'b1;
		10'd292: fft_load[36] = 1'b1;
		10'd293: fft_load[37] = 1'b1;
		10'd294: fft_load[38] = 1'b1;
		10'd295: fft_load[39] = 1'b1;
		10'd296: fft_load[40] = 1'b1;
		10'd297: fft_load[41] = 1'b1;
		10'd298: fft_load[42] = 1'b1;
		10'd299: fft_load[43] = 1'b1;
		10'd300: fft_load[44] = 1'b1;
		10'd301: fft_load[45] = 1'b1;
		10'd302: fft_load[46] = 1'b1;
		10'd303: fft_load[47] = 1'b1;
		10'd304: fft_load[48] = 1'b1;
		10'd305: fft_load[49] = 1'b1;
		10'd306: fft_load[50] = 1'b1;
		10'd307: fft_load[51] = 1'b1;
		10'd308: fft_load[52] = 1'b1;
		10'd309: fft_load[53] = 1'b1;
		10'd310: fft_load[54] = 1'b1;
		10'd311: fft_load[55] = 1'b1;
		10'd312: fft_load[56] = 1'b1;
		10'd313: fft_load[57] = 1'b1;
		10'd314: fft_load[58] = 1'b1;
		10'd315: fft_load[59] = 1'b1;
		10'd316: fft_load[60] = 1'b1;
		10'd317: fft_load[61] = 1'b1;
		10'd318: fft_load[62] = 1'b1;
		10'd319: fft_load[63] = 1'b1;
		10'd320: fft_load[64] = 1'b1;
		10'd321: fft_load[65] = 1'b1;
		10'd322: fft_load[66] = 1'b1;
		10'd323: fft_load[67] = 1'b1;
		10'd324: fft_load[68] = 1'b1;
		10'd325: fft_load[69] = 1'b1;
		10'd326: fft_load[70] = 1'b1;
		10'd327: fft_load[71] = 1'b1;
		10'd328: fft_load[72] = 1'b1;
		10'd329: fft_load[73] = 1'b1;
		10'd330: fft_load[74] = 1'b1;
		10'd331: fft_load[75] = 1'b1;
		10'd332: fft_load[76] = 1'b1;
		10'd333: fft_load[77] = 1'b1;
		10'd334: fft_load[78] = 1'b1;
		10'd335: fft_load[79] = 1'b1;
		10'd336: fft_load[80] = 1'b1;
		10'd337: fft_load[81] = 1'b1;
		10'd338: fft_load[82] = 1'b1;
		10'd339: fft_load[83] = 1'b1;
		10'd340: fft_load[84] = 1'b1;
		10'd341: fft_load[85] = 1'b1;
		10'd342: fft_load[86] = 1'b1;
		10'd343: fft_load[87] = 1'b1;
		10'd344: fft_load[88] = 1'b1;
		10'd345: fft_load[89] = 1'b1;
		10'd346: fft_load[90] = 1'b1;
		10'd347: fft_load[91] = 1'b1;
		10'd348: fft_load[92] = 1'b1;
		10'd349: fft_load[93] = 1'b1;
		10'd350: fft_load[94] = 1'b1;
		10'd351: fft_load[95] = 1'b1;
		10'd352: fft_load[96] = 1'b1;
		10'd353: fft_load[97] = 1'b1;
		10'd354: fft_load[98] = 1'b1;
		10'd355: fft_load[99] = 1'b1;
		10'd356: fft_load[100] = 1'b1;
		10'd357: fft_load[101] = 1'b1;
		10'd358: fft_load[102] = 1'b1;
		10'd359: fft_load[103] = 1'b1;
		10'd360: fft_load[104] = 1'b1;
		10'd361: fft_load[105] = 1'b1;
		10'd362: fft_load[106] = 1'b1;
		10'd363: fft_load[107] = 1'b1;
		10'd364: fft_load[108] = 1'b1;
		10'd365: fft_load[109] = 1'b1;
		10'd366: fft_load[110] = 1'b1;
		10'd367: fft_load[111] = 1'b1;
		10'd368: fft_load[112] = 1'b1;
		10'd369: fft_load[113] = 1'b1;
		10'd370: fft_load[114] = 1'b1;
		10'd371: fft_load[115] = 1'b1;
		10'd372: fft_load[116] = 1'b1;
		10'd373: fft_load[117] = 1'b1;
		10'd374: fft_load[118] = 1'b1;
		10'd375: fft_load[119] = 1'b1;
		10'd376: fft_load[120] = 1'b1;
		10'd377: fft_load[121] = 1'b1;
		10'd378: fft_load[122] = 1'b1;
		10'd379: fft_load[123] = 1'b1;
		10'd380: fft_load[124] = 1'b1;
		10'd381: fft_load[125] = 1'b1;
		10'd382: fft_load[126] = 1'b1;
		10'd383: fft_load[127] = 1'b1;
		10'd384: fft_load[128] = 1'b1;
		10'd385: fft_load[129] = 1'b1;
		10'd386: fft_load[130] = 1'b1;
		10'd387: fft_load[131] = 1'b1;
		10'd388: fft_load[132] = 1'b1;
		10'd389: fft_load[133] = 1'b1;
		10'd390: fft_load[134] = 1'b1;
		10'd391: fft_load[135] = 1'b1;
		10'd392: fft_load[136] = 1'b1;
		10'd393: fft_load[137] = 1'b1;
		10'd394: fft_load[138] = 1'b1;
		10'd395: fft_load[139] = 1'b1;
		10'd396: fft_load[140] = 1'b1;
		10'd397: fft_load[141] = 1'b1;
		10'd398: fft_load[142] = 1'b1;
		10'd399: fft_load[143] = 1'b1;
		10'd400: fft_load[144] = 1'b1;
		10'd401: fft_load[145] = 1'b1;
		10'd402: fft_load[146] = 1'b1;
		10'd403: fft_load[147] = 1'b1;
		10'd404: fft_load[148] = 1'b1;
		10'd405: fft_load[149] = 1'b1;
		10'd406: fft_load[150] = 1'b1;
		10'd407: fft_load[151] = 1'b1;
		10'd408: fft_load[152] = 1'b1;
		10'd409: fft_load[153] = 1'b1;
		10'd410: fft_load[154] = 1'b1;
		10'd411: fft_load[155] = 1'b1;
		10'd412: fft_load[156] = 1'b1;
		10'd413: fft_load[157] = 1'b1;
		10'd414: fft_load[158] = 1'b1;
		10'd415: fft_load[159] = 1'b1;
		10'd416: fft_load[160] = 1'b1;
		10'd417: fft_load[161] = 1'b1;
		10'd418: fft_load[162] = 1'b1;
		10'd419: fft_load[163] = 1'b1;
		10'd420: fft_load[164] = 1'b1;
		10'd421: fft_load[165] = 1'b1;
		10'd422: fft_load[166] = 1'b1;
		10'd423: fft_load[167] = 1'b1;
		10'd424: fft_load[168] = 1'b1;
		10'd425: fft_load[169] = 1'b1;
		10'd426: fft_load[170] = 1'b1;
		10'd427: fft_load[171] = 1'b1;
		10'd428: fft_load[172] = 1'b1;
		10'd429: fft_load[173] = 1'b1;
		10'd430: fft_load[174] = 1'b1;
		10'd431: fft_load[175] = 1'b1;
		10'd432: fft_load[176] = 1'b1;
		10'd433: fft_load[177] = 1'b1;
		10'd434: fft_load[178] = 1'b1;
		10'd435: fft_load[179] = 1'b1;
		10'd436: fft_load[180] = 1'b1;
		10'd437: fft_load[181] = 1'b1;
		10'd438: fft_load[182] = 1'b1;
		10'd439: fft_load[183] = 1'b1;
		10'd440: fft_load[184] = 1'b1;
		10'd441: fft_load[185] = 1'b1;
		10'd442: fft_load[186] = 1'b1;
		10'd443: fft_load[187] = 1'b1;
		10'd444: fft_load[188] = 1'b1;
		10'd445: fft_load[189] = 1'b1;
		10'd446: fft_load[190] = 1'b1;
		10'd447: fft_load[191] = 1'b1;
		10'd448: fft_load[192] = 1'b1;
		10'd449: fft_load[193] = 1'b1;
		10'd450: fft_load[194] = 1'b1;
		10'd451: fft_load[195] = 1'b1;
		10'd452: fft_load[196] = 1'b1;
		10'd453: fft_load[197] = 1'b1;
		10'd454: fft_load[198] = 1'b1;
		10'd455: fft_load[199] = 1'b1;
		10'd456: fft_load[200] = 1'b1;
		10'd457: fft_load[201] = 1'b1;
		10'd458: fft_load[202] = 1'b1;
		10'd459: fft_load[203] = 1'b1;
		10'd460: fft_load[204] = 1'b1;
		10'd461: fft_load[205] = 1'b1;
		10'd462: fft_load[206] = 1'b1;
		10'd463: fft_load[207] = 1'b1;
		10'd464: fft_load[208] = 1'b1;
		10'd465: fft_load[209] = 1'b1;
		10'd466: fft_load[210] = 1'b1;
		10'd467: fft_load[211] = 1'b1;
		10'd468: fft_load[212] = 1'b1;
		10'd469: fft_load[213] = 1'b1;
		10'd470: fft_load[214] = 1'b1;
		10'd471: fft_load[215] = 1'b1;
		10'd472: fft_load[216] = 1'b1;
		10'd473: fft_load[217] = 1'b1;
		10'd474: fft_load[218] = 1'b1;
		10'd475: fft_load[219] = 1'b1;
		10'd476: fft_load[220] = 1'b1;
		10'd477: fft_load[221] = 1'b1;
		10'd478: fft_load[222] = 1'b1;
		10'd479: fft_load[223] = 1'b1;
		10'd480: fft_load[224] = 1'b1;
		10'd481: fft_load[225] = 1'b1;
		10'd482: fft_load[226] = 1'b1;
		10'd483: fft_load[227] = 1'b1;
		10'd484: fft_load[228] = 1'b1;
		10'd485: fft_load[229] = 1'b1;
		10'd486: fft_load[230] = 1'b1;
		10'd487: fft_load[231] = 1'b1;
		10'd488: fft_load[232] = 1'b1;
		10'd489: fft_load[233] = 1'b1;
		10'd490: fft_load[234] = 1'b1;
		10'd491: fft_load[235] = 1'b1;
		10'd492: fft_load[236] = 1'b1;
		10'd493: fft_load[237] = 1'b1;
		10'd494: fft_load[238] = 1'b1;
		10'd495: fft_load[239] = 1'b1;
		10'd496: fft_load[240] = 1'b1;
		10'd497: fft_load[241] = 1'b1;
		10'd498: fft_load[242] = 1'b1;
		10'd499: fft_load[243] = 1'b1;
		10'd500: fft_load[244] = 1'b1;
		10'd501: fft_load[245] = 1'b1;
		10'd502: fft_load[246] = 1'b1;
		10'd503: fft_load[247] = 1'b1;
		10'd504: fft_load[248] = 1'b1;
		10'd505: fft_load[249] = 1'b1;
		10'd506: fft_load[250] = 1'b1;
		10'd507: fft_load[251] = 1'b1;
		10'd508: fft_load[252] = 1'b1;
		10'd509: fft_load[253] = 1'b1;
		10'd510: fft_load[254] = 1'b1;
		10'd511: fft_load[255] = 1'b1;
		default: ;
	endcase
	case (AVL_ADDR)
		10'd512: READY_load = 1'b1;
		default: READY_load = 1'b0;
	endcase

end
endmodule
